`timescale 1ns / 1ps
module tb_parity_generator;

reg in0, in1, in2;
wire parity_out;

parity_generator dut (
    .in0(in0),
    .in1(in1),
    .in2(in2),
    .parity_out(parity_out)
);

initial begin
    // Test cases
    in0 = 0; in1 = 0; in2 = 0; #10;
    in0 = 0; in1 = 0; in2 = 1; #10;
    in0 = 1; in1 = 1; in2 = 0; #10;
    in0 = 1; in1 = 1; in2 = 1; #10;
    $finish;
end

endmodule
